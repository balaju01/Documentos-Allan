LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY CONTADOR_D IS
	GENERIC( N : INTEGER := 4 );
	PORT(
		EN,CLR,CLK: IN STD_LOGIC;
		DISPLAY : INOUT STD_LOGIC_VECTOR(8 DOWNTO 0)
	);
END CONTADOR_D;

ARCHITECTURE PROGRAMA OF CONTADOR_A IS
CONSTANT A : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0001000";
CONSTANT L : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "1001111";
CONSTANT N : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "1101010";
CONSTANT Z : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0010010";
CONSTANT E : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0110000";
CONSTANT P : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0011000";
CONSTANT D : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "1000010";
CONSTANT E1 : STD_LOGIC_VECTOR( 1 DOWNTO 0 ) := "00";
CONSTANT E2 : STD_LOGIC_VECTOR( 1 DOWNTO 0 ) := "01";
CONSTANT E3 : STD_LOGIC_VECTOR( 1 DOWNTO 0 ) := "10";
CONSTANT ERROR : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "11111111";
CONSTANT D0 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := E1&A;
CONSTANT D1 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := E1&L;
CONSTANT D2 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := E2&L;
CONSTANT D3 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := E2&A;
CONSTANT D4 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := E1&N;
CONSTANT D5 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := E1&Z;
CONSTANT D6 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := E1&E;
CONSTANT D7 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := E1&P;
CONSTANT D8 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := E2&E;
CONSTANT D9 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := E1&D;
CONSTANT D10 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := E3&A;
BEGIN
	PCONT_D : PROCESS( CLK, CLR )
	BEGIN
		IF( CLR = '1' )THEN
			DISPLAY <= D0;
		ELSIF( CLK'EVENT AND CLK = '1' )THEN
			IF( EN = '1' )THEN			
				CASE DISPLAY IS
					WHEN D0 =>
							DISPLAY <= D1
					WHEN D1 =>
							DISPLAY <= D2
					WHEN D2 =>
							DISPLAY <= D3
					WHEN D3 =>
							DISPLAY <= D4
					WHEN D4 =>
							DISPLAY <= D5
					WHEN D5 =>
							DISPLAY <= D6
					WHEN D6 =>
							DISPLAY <= D7
					WHEN D7 =>
							DISPLAY <= D8
					WHEN D8 =>
							DISPLAY <= D9
					WHEN D9 =>
							DISPLAY <= D10
					WHEN D10 =>
							DISPLAY <= D0
					WHEN OTHERS=>
						--	DISPLAY <= "-------";
							DISPLAY <= D0;
						--	DISPLAY <= ERROR;
				END CASE;
			END IF;
		END IF;
	END PROCESS PCONT_D;
END PROGRAMA;