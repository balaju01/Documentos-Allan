LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY CONTADOR_E IS
	GENERIC( N : INTEGER := 4 );
	PORT(
		EN,CLR,CLK: IN STD_LOGIC;
		DISPLAY : INOUT STD_LOGIC_VECTOR(8 DOWNTO 0)
	);
END CONTADOR_E;

ARCHITECTURE PROGRAMA OF CONTADOR_A IS
CONSTANT S2 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0010010";
CONSTANT S0 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0000001";
CONSTANT S1 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "1001111";
CONSTANT S6 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0100000";
CONSTANT S3 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0000110";
CONSTANT S5 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0100100";
CONSTANT S8 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0000000";
CONSTANT E1 : STD_LOGIC_VECTOR( 1 DOWNTO 0 ) := "00";
CONSTANT E2 : STD_LOGIC_VECTOR( 1 DOWNTO 0 ) := "01";
CONSTANT E3 : STD_LOGIC_VECTOR( 1 DOWNTO 0 ) := "10";
CONSTANT ERROR : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "11111111";
CONSTANT D0 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := E1&S2;
CONSTANT D1 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := E1&S0;
CONSTANT D2 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := E1&S1;
CONSTANT D3 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := E2&S1;
CONSTANT D4 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := E1&S6;
CONSTANT D5 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := E1&S3;
CONSTANT D6 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := E2&S0;
CONSTANT D7 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := E1&S5;
CONSTANT D8 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := E1&S8;
CONSTANT D9 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := E2&S8;

BEGIN
	PCONT_E : PROCESS( CLK, CLR )
	BEGIN
		IF( CLR = '1' )THEN
			DISPLAY <= D0;
		ELSIF( CLK'EVENT AND CLK = '1' )THEN
			IF( EN = '1' )THEN			
				CASE DISPLAY IS
					WHEN D0 =>
							DISPLAY <= D1
					WHEN D1 =>
							DISPLAY <= D2
					WHEN D2 =>
							DISPLAY <= D3
					WHEN D3 =>
							DISPLAY <= D4
					WHEN D4 =>
							DISPLAY <= D5
					WHEN D5 =>
							DISPLAY <= D6
					WHEN D6 =>
							DISPLAY <= D7
					WHEN D7 =>
							DISPLAY <= D8
					WHEN D8 =>
							DISPLAY <= D9
					WHEN D9 =>
							DISPLAY <= D0
					
					WHEN OTHERS=>
						--	DISPLAY <= "-------";
							DISPLAY <= D0;
						--	DISPLAY <= ERROR;
				END CASE;
			END IF;
		END IF;
	END PROCESS PCONT_E;
END PROGRAMA;