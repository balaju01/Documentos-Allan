library ieee;
use ieee.std_logic_1164.all;

entity mensaje is
	port(
		CLK,CLR IN STD_LOGIC;
		AN OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		DISP OUT STD_LOGIC_VECTOR (6 DOWNTO 0)
	);
end mensaje;

ARCHITECTURE PROGRAMA OF MENSAJE IS
--CONSTANT LETRA_N:STD_LOGIC_VECTOR(6 DOWNTO 0):="
BEGIN
	IPN:PROCESS(CLR,CLK)
	BEGIN
		IF (CLR='1') THEN
			AN<="110";
		ELSIF(CLK'EVENT AND CLK='1')THEN
			AN(0)<=AN(3);
			AN(1)<=AN(0);
			AN(2)<=AN(1);
			AN(3)<=AN(2);
		END IF;
	END PROCESS IPN;
	DISP<="1101010" WHEN (AN="101") ELSE
			"0011000"WHEN (AN="011") ELSE
			"1001111"WHEN (AN="110") ELSE
			"0000000"
END PROGRAMA;