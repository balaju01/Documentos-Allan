LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY CONTADOR_C IS
	GENERIC( N : INTEGER := 4 );
	PORT(
		EN,CLR,CLK: IN STD_LOGIC;
		DISPLAY : INOUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END CONTADOR_C;

ARCHITECTURE PROGRAMA OF CONTADOR_C IS
CONSTANT D0 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "1001111";
CONSTANT D1 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0010010";
CONSTANT D2 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0000110";
CONSTANT D3 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "1001100";
CONSTANT D4 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0100100";
CONSTANT D5 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0100000";

CONSTANT ERROR : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "11111111";

BEGIN
	PCONT_C : PROCESS( CLK, CLR )
	BEGIN
		IF( CLR = '1' )THEN
			DISPLAY <= D0;
		ELSIF( CLK'EVENT AND CLK = '1' )THEN
			IF( EN = '1' )THEN			
				CASE DISPLAY IS
					WHEN D0 =>
							DISPLAY <= D1
					WHEN D1 =>
							DISPLAY <= D2
					WHEN D2 =>
							DISPLAY <= D3
					WHEN D3 =>
							DISPLAY <= D4
					WHEN D4 =>
							DISPLAY <= D5
					WHEN D5 =>
							DISPLAY <= D0
					WHEN OTHERS=>
						--	DISPLAY <= "-------";
							DISPLAY <= D0;
						--	DISPLAY <= ERROR;
				END CASE;
			END IF;
		END IF;
	END PROCESS PCONT_C;
END PROGRAMA;