LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY CONTADOR IS
	GENERIC( N : INTEGER := 4 );
	PORT(
		EN,CLR,CLK: IN STD_LOGIC;
		DISPLAY : INOUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END CONTADOR;

ARCHITECTURE PROGRAMA OF CONTADOR IS
CONSTANT D0 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0000001";
CONSTANT D1 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "1001111";
CONSTANT D2 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0010010";
CONSTANT D3 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0000110";
CONSTANT D4 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "1001100";
CONSTANT D5 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0100100";
CONSTANT D6 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0100000";
CONSTANT D7 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0001111";
CONSTANT D8 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0000000";
CONSTANT D9 : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0001100";
CONSTANT DA : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0001000";
CONSTANT DB : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "1100000";
CONSTANT DC : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "1100001";
CONSTANT DD : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "1000010";
CONSTANT DE : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0110000";
CONSTANT DF : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0111000";
CONSTANT ERROR : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "11111111";

BEGIN
	PCONT : PROCESS( CLK, CLR )
	BEGIN
		IF( CLR = '1' )THEN
			DISPLAY <= D0;
		ELSIF( CLK'EVENT AND CLK = '1' )THEN
			IF( EN = '1' )THEN			
				CASE DISPLAY IS
					WHEN D0 =>
							DISPLAY <= D1
					WHEN D1 =>
							DISPLAY <= D2
					WHEN D2 =>
							DISPLAY <= D3
							--CONTINUARA...
					WHEN OTHERS=>
						--	DISPLAY <= "-------";
							DISPLAY <= D0;
						--	DISPLAY <= ERROR;
				END CASE;
			END IF;
		END IF;
	END PROCESS PCONT;
END PROGRAMA;