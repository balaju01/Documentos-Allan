LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY MARQUESINA IS
	PORT(CLK, CLR : IN STD_LOGIC;
	E: IN STD_LOGIC_VECTOR (2 DOWN TO 0);
	SAL : OUT STD_LOGIC_VECTOR(9 DOWN TO 0);
	AN OUT STD_LOGIC_VECTOR (2 DOWNTO 0)
	);
END MARQUESINA;

ARCHITECTURE CONTADOR OF BOLETA IS
CONSTANT LETRA_H: STD_LOGIC_VECTOR(6 DOWNTO 0):="1001000";
CONSTANT LETRA_0: STD_LOGIC_VECTOR(6 DOWNTO 0):="0000001";
CONSTANT LETRA_L: STD_LOGIC_VECTOR(6 DOWNTO 0):="1110001";
CONSTANT LETRA_A: STD_LOGIC_VECTOR(6 DOWNTO 0):="0001000";
CONSTANT NL: STD_LOGIC_VECTOR(6 DOWNTO 0):="1111111";

CONSTANT D0: STD_LOGIC_VECTOR(2 DOWNTO 0):="110";
CONSTANT D1: STD_LOGIC_VECTOR(2 DOWNTO 0):="101";
CONSTANT D2: STD_LOGIC_VECTOR(2 DOWNTO 0):="011";
CONSTANT ND: STD_LOGIC_VECTOR(2 DOWNTO 0):="111";

CONSTANT Q0: STD_LOGIC_VECTOR(9 DOWNTO 0):=ND&NL;
CONSTANT Q1: STD_LOGIC_VECTOR(9 DOWNTO 0):=D0&LETRA_H;
CONSTANT Q2: STD_LOGIC_VECTOR(9 DOWNTO 0):=D1&LETRA_H;
CONSTANT Q3: STD_LOGIC_VECTOR(9 DOWNTO 0):=D0&LETRA_0;
CONSTANT Q4: STD_LOGIC_VECTOR(9 DOWNTO 0):=D2&LETRA_H;
CONSTANT Q5: STD_LOGIC_VECTOR(9 DOWNTO 0):=D1&LETRA_0;
CONSTANT Q6: STD_LOGIC_VECTOR(9 DOWNTO 0):=D0&LETRA_L;
CONSTANT Q7: STD_LOGIC_VECTOR(9 DOWNTO 0):=D2&LETRA_0;
CONSTANT Q8: STD_LOGIC_VECTOR(9 DOWNTO 0):=D1&LETRA_L;
CONSTANT Q9: STD_LOGIC_VECTOR(9 DOWNTO 0):=D0&LETRA_A;
CONSTANT Q10: STD_LOGIC_VECTOR(9 DOWNTO 0):=D2&LETRA_L;
CONSTANT Q11: STD_LOGIC_VECTOR(9 DOWNTO 0):=D1&LETRA_A;
CONSTANT Q12: STD_LOGIC_VECTOR(9 DOWNTO 0):=D2&LETRA_A;

002180700816243897
002180700816243897

BEGIN
	CONT:PROCES(CLK,CLR)
	BEGIN
		IF(CLR='1')THEN
			SAL<=Q0;
		ELSIF(CLK'EVENT AND CLK='1')THEN
			CASE SAL IS
				WHEN Q0=>
					IF(E="000" OR E="001")THEN
						SAL<=Q0;
						AN<="111";
					ELSIF(E="010")THEN
						SAL<=Q1;
					ELSE
						SAL<=Q0;
					END IF;
				WHEN Q1=>
					IF(E="011")THEN
						SAL <= Q2;
					ELSIF(E="010")THEN
						SAL <= Q1;
					ELSE
						SAL <= Q1;
					END IF;
				WHEN Q2=>
					IF(E<="100")THEN
						SAL<=Q4;
					ELSIF(E<="011")THEN
						SAL<=Q3;
					ELSE
						SAL<=Q3;
					END IF;
				WHEN Q3=>
					IF(E<="100")THEN
						SAL<=Q4;
					ELSIF(E<="011")THEN
						SAL<=Q2;
					ELSE
						SAL<=Q2;
					END IF;
				WHEN Q4=>
					IF(E<="101")THEN
						SAL<=Q7;
					ELSIF(E<="100")THEN
						SAL<=Q5;
					ELSE
						SAL<=Q5;
					END IF;
				WHEN Q5=>
					IF(E<="101")THEN
						SAL<=Q7;
					ELSIF(E<="100")THEN
						SAL<=Q6;
					ELSE
						SAL<=Q6;
					END IF;
				WHEN Q6=>
					IF(E<="101")THEN
						SAL<=Q7;
					ELSIF(E<="100")THEN
						SAL<=Q4;
					ELSE
						SAL<=Q4;
					END IF;
				WHEN Q7=>
					IF(E<="110")THEN
						SAL<=Q10;
					ELSIF(E<="101")THEN
						SAL<=Q8;
					ELSE
						SAL<=Q8;
					END IF;
				WHEN Q8=>
					IF(E<="110")THEN
						SAL<=Q10;
					ELSIF(E<="101")THEN
						SAL<=Q9;
					ELSE
						SAL<=Q9;
					END IF;
				WHEN Q9=>
					IF(E<="110")THEN
						SAL<=Q10;
					ELSIF(E<="101")THEN
						SAL<=Q7;
					ELSE
						SAL<=Q7;
					END IF;
				WHEN Q10=>
					IF(E<="111")THEN
						SAL<=Q12;
					ELSIF(E<="110")THEN
						SAL<=Q11;
					ELSE
						SAL<=Q11;
					END IF;
				WHEN Q11=>
					IF(E<="111")THEN
						SAL<=Q12;
					ELSIF(E<="110")THEN
						SAL<=Q10;
					ELSE
						SAL<=Q10;
					END IF;
				WHEN Q12=>
					IF(E<="111")THEN
						SAL<=Q12;
					ELSIF(E<="000")THEN
						SAL<=Q0;
					ELSE
						SAL<=Q0;
					END IF;
				WHEN OTHERS=>
					SAL<=Q0;
			END CASE;	
		END IF;
	END PROCESS CONT;
	AS(2)<=SAL(9);
	AS(1)<=SAL(8);
	AS(0)<=SAL(7);
END CONTADOR;